library verilog;
use verilog.vl_types.all;
entity tb_single_cycle is
end tb_single_cycle;
