library verilog;
use verilog.vl_types.all;
entity single_cycle_tb is
end single_cycle_tb;
