library verilog;
use verilog.vl_types.all;
entity milestone1_test_vlg_vec_tst is
end milestone1_test_vlg_vec_tst;
