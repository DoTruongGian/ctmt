module single_cycle (

);


endmodule