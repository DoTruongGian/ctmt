library verilog;
use verilog.vl_types.all;
entity single_cycle_vlg_vec_tst is
end single_cycle_vlg_vec_tst;
