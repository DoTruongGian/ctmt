module convert7seg (
    input logic [6:0]  o_io_hex0,
    input logic [6:0]  o_io_hex1,
    input logic [6:0]  o_io_hex2,
    input logic [6:0]  o_io_hex3,
    input logic [6:0]  o_io_hex4,
    input logic [6:0]  o_io_hex5,
    input logic [6:0]  o_io_hex6,
    input logic [6:0]  o_io_hex7,
	 output logic [6:0]  o_io_hex0,
    output logic [6:0]  o_io_hex1,
    output logic [6:0]  o_io_hex2,
    output logic [6:0]  o_io_hex3,
    output logic [6:0]  o_io_hex4,
    output logic [6:0]  o_io_hex5,
    output logic [6:0]  o_io_hex6,
    output logic [6:0]  o_io_hex7
);

endmodule
